module lib

pub struct Generator {

}

pub fn (g Generator) generate(f FileParser) {
	//print(f)
	//exit(2)
}